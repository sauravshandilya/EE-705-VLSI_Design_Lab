-- Author: Saurav Shandilya
-- Description: mynor (NOR Gate implementation)


--import std_logic from the IEEE library
library ieee;
use ieee.std_logic_1164.all;

--ENTITY DECLARATION: name, inputs, outputs
entity mynor is					
   port( in1, in2 : in bit;
            out1 : out bit);
end mynor;

--Architecture of AND gate
architecture arch of mynor is 
begin
  out1 <= in1 nor in2;		
end arch;
