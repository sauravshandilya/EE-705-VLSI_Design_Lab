library verilog;
use verilog.vl_types.all;
entity helloworld is
end helloworld;
