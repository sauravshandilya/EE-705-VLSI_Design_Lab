-------------------------
-- Author: Saurav Shandilya
-- Description: BM Datapath implementation
-------------------------

-- ****** Datapath *******
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity bmdatapath is
      port ( 
	sysclk: In std_logic;		-- input to data block
	add:
	sub:

	---- Signal to controller	
	boothbit : In std_logic;
	qlsb: In std_logic;		

	---- Signal from controller
	       	
	     );
end bmdatapath;

architecture arch of bmdatapath is


	
end arch;
