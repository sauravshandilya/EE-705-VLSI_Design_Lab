-- Author: Saurav Shandilya
-- Description: myxor (XOR Gate implementation)


--import std_logic from the IEEE library
library ieee;
use ieee.std_logic_1164.all;

--ENTITY DECLARATION: name, inputs, outputs
entity myxor is					
   port( in1, in2 : in bit;
            out1 : out bit);
end myxor;

--Architecture of AND gate
architecture arch of myxor is 
begin
  out1 <= in1 xor in2;		
end arch;
