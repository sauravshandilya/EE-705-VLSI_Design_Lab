/*
-- Author: Saurav Shandilya 
-- Roll No: 153076004, Electronics System, EE, IIT Bombay
-- EE-705 VLSI Design Lab (Course Instructor: Prof. Virendra Singh)
-- Description: 6 FLoor Lift controller using verilog
--              System consist of 6 floor (Ground floor to 5th Floor).
--              
*/

module elevator6floor 
(
	reset,
	clk,
	carcall,
	hallcall_up,
	hallcall_down,
	floorsensor,

	carled,
	hallcall_upled,
	hallcall_downled,
	floorindicatorled,
	dooropen,
	dir_up,
	dir_down,
	liftmoving
);

endmodule



