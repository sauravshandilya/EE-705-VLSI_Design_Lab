---
-- Author: Saurav Shandilya
-- Description: Converts negative number into positive number. Negative number is detected by MSB bit
--              of register. If number is negative, perform two's complement. Mux either output 
--              2's complement (for -ve number) or nmber itself (for +ve number)
  


---

---library 
Library ieee;
USE IEEE.STD_LOGIC_1164.ALL;

--- entity

entity toPositive is
port 
(
    input : in bit_vector(7 downto 0);
    isnegative : out bit;
    output : out bit_vector(7 downto 0);
    clk : in bit;
    reset : in bit;   
    enable : in bit  
);
end toPositive;

architecture arch of toPositive is


component reg 
    generic ( nbits : integer); 
     port (
    data_in : in bit_vector(nbits-1 downto 0);
    data_out : out bit_vector(nbits-1 downto 0);
    clk : in bit;
    enable : in  bit;
    reset : in  bit
    );
  end component;

component mynot is					
   port( in1 : in bit;
        out1 : out bit);
end component;

component fullAdder_8bit
   port( A, B : in bit_vector(7 downto 0);
         sum: out bit_vector(7 downto 0); 
	 Cout : out bit);
end component;

component Mux2x1_8bit is
	port 
	( Mux_in_1:IN bit_vector(7 DOWNTO 0);
		Mux_in_2:IN bit_vector(7 DOWNTO 0);
		sel:IN bit; 
		mux_out:OUT bit_vector(7 DOWNTO 0)
	);		
end component;

signal reg_dataout : bit_vector(7 downto 0);
signal not_8bitout : bit_vector(7 downto 0);
signal twocomp_out : bit_vector(7 downto 0);

begin
  
inputdata: reg
    generic map ( nbits => 8 )
    port map (
      data_in => input,     -- 8 MSB bits are zero
      data_out => reg_dataout,             
      clk      => clk,
      reset    => reset,
      enable   => enable);

-- 1's complement    
grp_gen: for i in 0 to 7 generate
		grp_mynot: mynot port map (reg_dataout(i),not_8bitout(i));
	end generate grp_gen;    

-- 2's complement
 twocomp: fullAdder_8bit port map(not_8bitout,"00000001", twocomp_out);
 
-- If number is Postive, out<=number; else out<= 2's complement(number)  
 mux1: Mux2x1_8bit port map (reg_dataout,twocomp_out,reg_dataout(7),output);   -- reg_dataout(7) 1<= -ve number
  
end arch;